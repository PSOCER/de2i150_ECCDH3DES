// $Id: mg78$
// Created: 3/18/2015
// Author: Nico Bellante
// Lab Section: 337-03
// Description: sbox substitutions


module des_sbox_substitutions (
    input logic [0:47] input_wires,
    output logic [0:31] output_wires
);

// applies sbox substitutions as per the standards set for DES
always_comb
begin
case(input_wires[0:5])
    6'b000000: output_wires[0:3] = 4'd14;
    6'b000001: output_wires[0:3] = 4'd0;
    6'b000010: output_wires[0:3] = 4'd4;
    6'b000011: output_wires[0:3] = 4'd15;
    6'b000100: output_wires[0:3] = 4'd13;
    6'b000101: output_wires[0:3] = 4'd7;
    6'b000110: output_wires[0:3] = 4'd1;
    6'b000111: output_wires[0:3] = 4'd4;
    6'b001000: output_wires[0:3] = 4'd2;
    6'b001001: output_wires[0:3] = 4'd14;
    6'b001010: output_wires[0:3] = 4'd15;
    6'b001011: output_wires[0:3] = 4'd2;
    6'b001100: output_wires[0:3] = 4'd11;
    6'b001101: output_wires[0:3] = 4'd13;
    6'b001110: output_wires[0:3] = 4'd8;
    6'b001111: output_wires[0:3] = 4'd1;
    6'b010000: output_wires[0:3] = 4'd3;
    6'b010001: output_wires[0:3] = 4'd10;
    6'b010010: output_wires[0:3] = 4'd10;
    6'b010011: output_wires[0:3] = 4'd6;
    6'b010100: output_wires[0:3] = 4'd6;
    6'b010101: output_wires[0:3] = 4'd12;
    6'b010110: output_wires[0:3] = 4'd12;
    6'b010111: output_wires[0:3] = 4'd11;
    6'b011000: output_wires[0:3] = 4'd5;
    6'b011001: output_wires[0:3] = 4'd9;
    6'b011010: output_wires[0:3] = 4'd9;
    6'b011011: output_wires[0:3] = 4'd5;
    6'b011100: output_wires[0:3] = 4'd0;
    6'b011101: output_wires[0:3] = 4'd3;
    6'b011110: output_wires[0:3] = 4'd7;
    6'b011111: output_wires[0:3] = 4'd8;
    6'b100000: output_wires[0:3] = 4'd4;
    6'b100001: output_wires[0:3] = 4'd15;
    6'b100010: output_wires[0:3] = 4'd1;
    6'b100011: output_wires[0:3] = 4'd12;
    6'b100100: output_wires[0:3] = 4'd14;
    6'b100101: output_wires[0:3] = 4'd8;
    6'b100110: output_wires[0:3] = 4'd8;
    6'b100111: output_wires[0:3] = 4'd2;
    6'b101000: output_wires[0:3] = 4'd13;
    6'b101001: output_wires[0:3] = 4'd4;
    6'b101010: output_wires[0:3] = 4'd6;
    6'b101011: output_wires[0:3] = 4'd9;
    6'b101100: output_wires[0:3] = 4'd2;
    6'b101101: output_wires[0:3] = 4'd1;
    6'b101110: output_wires[0:3] = 4'd11;
    6'b101111: output_wires[0:3] = 4'd7;
    6'b110000: output_wires[0:3] = 4'd15;
    6'b110001: output_wires[0:3] = 4'd5;
    6'b110010: output_wires[0:3] = 4'd12;
    6'b110011: output_wires[0:3] = 4'd11;
    6'b110100: output_wires[0:3] = 4'd9;
    6'b110101: output_wires[0:3] = 4'd3;
    6'b110110: output_wires[0:3] = 4'd7;
    6'b110111: output_wires[0:3] = 4'd14;
    6'b111000: output_wires[0:3] = 4'd3;
    6'b111001: output_wires[0:3] = 4'd10;
    6'b111010: output_wires[0:3] = 4'd10;
    6'b111011: output_wires[0:3] = 4'd0;
    6'b111100: output_wires[0:3] = 4'd5;
    6'b111101: output_wires[0:3] = 4'd6;
    6'b111110: output_wires[0:3] = 4'd0;
    6'b111111: output_wires[0:3] = 4'd13;
endcase

case(input_wires[6:11])
    6'b000000: output_wires[4:7] = 4'd15;
    6'b000001: output_wires[4:7] = 4'd3;
    6'b000010: output_wires[4:7] = 4'd1;
    6'b000011: output_wires[4:7] = 4'd13;
    6'b000100: output_wires[4:7] = 4'd8;
    6'b000101: output_wires[4:7] = 4'd4;
    6'b000110: output_wires[4:7] = 4'd14;
    6'b000111: output_wires[4:7] = 4'd7;
    6'b001000: output_wires[4:7] = 4'd6;
    6'b001001: output_wires[4:7] = 4'd15;
    6'b001010: output_wires[4:7] = 4'd11;
    6'b001011: output_wires[4:7] = 4'd2;
    6'b001100: output_wires[4:7] = 4'd3;
    6'b001101: output_wires[4:7] = 4'd8;
    6'b001110: output_wires[4:7] = 4'd4;
    6'b001111: output_wires[4:7] = 4'd14;
    6'b010000: output_wires[4:7] = 4'd9;
    6'b010001: output_wires[4:7] = 4'd12;
    6'b010010: output_wires[4:7] = 4'd7;
    6'b010011: output_wires[4:7] = 4'd0;
    6'b010100: output_wires[4:7] = 4'd2;
    6'b010101: output_wires[4:7] = 4'd1;
    6'b010110: output_wires[4:7] = 4'd13;
    6'b010111: output_wires[4:7] = 4'd10;
    6'b011000: output_wires[4:7] = 4'd12;
    6'b011001: output_wires[4:7] = 4'd6;
    6'b011010: output_wires[4:7] = 4'd0;
    6'b011011: output_wires[4:7] = 4'd9;
    6'b011100: output_wires[4:7] = 4'd5;
    6'b011101: output_wires[4:7] = 4'd11;
    6'b011110: output_wires[4:7] = 4'd10;
    6'b011111: output_wires[4:7] = 4'd5;
    6'b100000: output_wires[4:7] = 4'd0;
    6'b100001: output_wires[4:7] = 4'd13;
    6'b100010: output_wires[4:7] = 4'd14;
    6'b100011: output_wires[4:7] = 4'd8;
    6'b100100: output_wires[4:7] = 4'd7;
    6'b100101: output_wires[4:7] = 4'd10;
    6'b100110: output_wires[4:7] = 4'd11;
    6'b100111: output_wires[4:7] = 4'd1;
    6'b101000: output_wires[4:7] = 4'd10;
    6'b101001: output_wires[4:7] = 4'd3;
    6'b101010: output_wires[4:7] = 4'd4;
    6'b101011: output_wires[4:7] = 4'd15;
    6'b101100: output_wires[4:7] = 4'd13;
    6'b101101: output_wires[4:7] = 4'd4;
    6'b101110: output_wires[4:7] = 4'd1;
    6'b101111: output_wires[4:7] = 4'd2;
    6'b110000: output_wires[4:7] = 4'd5;
    6'b110001: output_wires[4:7] = 4'd11;
    6'b110010: output_wires[4:7] = 4'd8;
    6'b110011: output_wires[4:7] = 4'd6;
    6'b110100: output_wires[4:7] = 4'd12;
    6'b110101: output_wires[4:7] = 4'd7;
    6'b110110: output_wires[4:7] = 4'd6;
    6'b110111: output_wires[4:7] = 4'd12;
    6'b111000: output_wires[4:7] = 4'd9;
    6'b111001: output_wires[4:7] = 4'd0;
    6'b111010: output_wires[4:7] = 4'd3;
    6'b111011: output_wires[4:7] = 4'd5;
    6'b111100: output_wires[4:7] = 4'd2;
    6'b111101: output_wires[4:7] = 4'd14;
    6'b111110: output_wires[4:7] = 4'd15;
    6'b111111: output_wires[4:7] = 4'd9;
endcase

case(input_wires[12:17])
    6'b000000: output_wires[8:11] = 4'd10;
    6'b000001: output_wires[8:11] = 4'd13;
    6'b000010: output_wires[8:11] = 4'd0;
    6'b000011: output_wires[8:11] = 4'd7;
    6'b000100: output_wires[8:11] = 4'd9;
    6'b000101: output_wires[8:11] = 4'd0;
    6'b000110: output_wires[8:11] = 4'd14;
    6'b000111: output_wires[8:11] = 4'd9;
    6'b001000: output_wires[8:11] = 4'd6;
    6'b001001: output_wires[8:11] = 4'd3;
    6'b001010: output_wires[8:11] = 4'd3;
    6'b001011: output_wires[8:11] = 4'd4;
    6'b001100: output_wires[8:11] = 4'd15;
    6'b001101: output_wires[8:11] = 4'd6;
    6'b001110: output_wires[8:11] = 4'd5;
    6'b001111: output_wires[8:11] = 4'd10;
    6'b010000: output_wires[8:11] = 4'd1;
    6'b010001: output_wires[8:11] = 4'd2;
    6'b010010: output_wires[8:11] = 4'd13;
    6'b010011: output_wires[8:11] = 4'd8;
    6'b010100: output_wires[8:11] = 4'd12;
    6'b010101: output_wires[8:11] = 4'd5;
    6'b010110: output_wires[8:11] = 4'd7;
    6'b010111: output_wires[8:11] = 4'd14;
    6'b011000: output_wires[8:11] = 4'd11;
    6'b011001: output_wires[8:11] = 4'd12;
    6'b011010: output_wires[8:11] = 4'd4;
    6'b011011: output_wires[8:11] = 4'd11;
    6'b011100: output_wires[8:11] = 4'd2;
    6'b011101: output_wires[8:11] = 4'd15;
    6'b011110: output_wires[8:11] = 4'd8;
    6'b011111: output_wires[8:11] = 4'd1;
    6'b100000: output_wires[8:11] = 4'd13;
    6'b100001: output_wires[8:11] = 4'd1;
    6'b100010: output_wires[8:11] = 4'd6;
    6'b100011: output_wires[8:11] = 4'd10;
    6'b100100: output_wires[8:11] = 4'd4;
    6'b100101: output_wires[8:11] = 4'd13;
    6'b100110: output_wires[8:11] = 4'd9;
    6'b100111: output_wires[8:11] = 4'd0;
    6'b101000: output_wires[8:11] = 4'd8;
    6'b101001: output_wires[8:11] = 4'd6;
    6'b101010: output_wires[8:11] = 4'd15;
    6'b101011: output_wires[8:11] = 4'd9;
    6'b101100: output_wires[8:11] = 4'd3;
    6'b101101: output_wires[8:11] = 4'd8;
    6'b101110: output_wires[8:11] = 4'd0;
    6'b101111: output_wires[8:11] = 4'd7;
    6'b110000: output_wires[8:11] = 4'd11;
    6'b110001: output_wires[8:11] = 4'd4;
    6'b110010: output_wires[8:11] = 4'd1;
    6'b110011: output_wires[8:11] = 4'd15;
    6'b110100: output_wires[8:11] = 4'd2;
    6'b110101: output_wires[8:11] = 4'd14;
    6'b110110: output_wires[8:11] = 4'd12;
    6'b110111: output_wires[8:11] = 4'd3;
    6'b111000: output_wires[8:11] = 4'd5;
    6'b111001: output_wires[8:11] = 4'd11;
    6'b111010: output_wires[8:11] = 4'd10;
    6'b111011: output_wires[8:11] = 4'd5;
    6'b111100: output_wires[8:11] = 4'd14;
    6'b111101: output_wires[8:11] = 4'd2;
    6'b111110: output_wires[8:11] = 4'd7;
    6'b111111: output_wires[8:11] = 4'd12;
endcase

case(input_wires[18:23])
    6'b000000: output_wires[12:15] = 4'd7;
    6'b000001: output_wires[12:15] = 4'd13;
    6'b000010: output_wires[12:15] = 4'd13;
    6'b000011: output_wires[12:15] = 4'd8;
    6'b000100: output_wires[12:15] = 4'd14;
    6'b000101: output_wires[12:15] = 4'd11;
    6'b000110: output_wires[12:15] = 4'd3;
    6'b000111: output_wires[12:15] = 4'd5;
    6'b001000: output_wires[12:15] = 4'd0;
    6'b001001: output_wires[12:15] = 4'd6;
    6'b001010: output_wires[12:15] = 4'd6;
    6'b001011: output_wires[12:15] = 4'd15;
    6'b001100: output_wires[12:15] = 4'd9;
    6'b001101: output_wires[12:15] = 4'd0;
    6'b001110: output_wires[12:15] = 4'd10;
    6'b001111: output_wires[12:15] = 4'd3;
    6'b010000: output_wires[12:15] = 4'd1;
    6'b010001: output_wires[12:15] = 4'd4;
    6'b010010: output_wires[12:15] = 4'd2;
    6'b010011: output_wires[12:15] = 4'd7;
    6'b010100: output_wires[12:15] = 4'd8;
    6'b010101: output_wires[12:15] = 4'd2;
    6'b010110: output_wires[12:15] = 4'd5;
    6'b010111: output_wires[12:15] = 4'd12;
    6'b011000: output_wires[12:15] = 4'd11;
    6'b011001: output_wires[12:15] = 4'd1;
    6'b011010: output_wires[12:15] = 4'd12;
    6'b011011: output_wires[12:15] = 4'd10;
    6'b011100: output_wires[12:15] = 4'd4;
    6'b011101: output_wires[12:15] = 4'd14;
    6'b011110: output_wires[12:15] = 4'd15;
    6'b011111: output_wires[12:15] = 4'd9;
    6'b100000: output_wires[12:15] = 4'd10;
    6'b100001: output_wires[12:15] = 4'd3;
    6'b100010: output_wires[12:15] = 4'd6;
    6'b100011: output_wires[12:15] = 4'd15;
    6'b100100: output_wires[12:15] = 4'd9;
    6'b100101: output_wires[12:15] = 4'd0;
    6'b100110: output_wires[12:15] = 4'd0;
    6'b100111: output_wires[12:15] = 4'd6;
    6'b101000: output_wires[12:15] = 4'd12;
    6'b101001: output_wires[12:15] = 4'd10;
    6'b101010: output_wires[12:15] = 4'd11;
    6'b101011: output_wires[12:15] = 4'd1;
    6'b101100: output_wires[12:15] = 4'd7;
    6'b101101: output_wires[12:15] = 4'd13;
    6'b101110: output_wires[12:15] = 4'd13;
    6'b101111: output_wires[12:15] = 4'd8;
    6'b110000: output_wires[12:15] = 4'd15;
    6'b110001: output_wires[12:15] = 4'd9;
    6'b110010: output_wires[12:15] = 4'd1;
    6'b110011: output_wires[12:15] = 4'd4;
    6'b110100: output_wires[12:15] = 4'd3;
    6'b110101: output_wires[12:15] = 4'd5;
    6'b110110: output_wires[12:15] = 4'd14;
    6'b110111: output_wires[12:15] = 4'd11;
    6'b111000: output_wires[12:15] = 4'd5;
    6'b111001: output_wires[12:15] = 4'd12;
    6'b111010: output_wires[12:15] = 4'd2;
    6'b111011: output_wires[12:15] = 4'd7;
    6'b111100: output_wires[12:15] = 4'd8;
    6'b111101: output_wires[12:15] = 4'd2;
    6'b111110: output_wires[12:15] = 4'd4;
    6'b111111: output_wires[12:15] = 4'd14;
endcase

case(input_wires[24:29])
    6'b000000: output_wires[16:19] = 4'd2;
    6'b000001: output_wires[16:19] = 4'd14;
    6'b000010: output_wires[16:19] = 4'd12;
    6'b000011: output_wires[16:19] = 4'd11;
    6'b000100: output_wires[16:19] = 4'd4;
    6'b000101: output_wires[16:19] = 4'd2;
    6'b000110: output_wires[16:19] = 4'd1;
    6'b000111: output_wires[16:19] = 4'd12;
    6'b001000: output_wires[16:19] = 4'd7;
    6'b001001: output_wires[16:19] = 4'd4;
    6'b001010: output_wires[16:19] = 4'd10;
    6'b001011: output_wires[16:19] = 4'd7;
    6'b001100: output_wires[16:19] = 4'd11;
    6'b001101: output_wires[16:19] = 4'd13;
    6'b001110: output_wires[16:19] = 4'd6;
    6'b001111: output_wires[16:19] = 4'd1;
    6'b010000: output_wires[16:19] = 4'd8;
    6'b010001: output_wires[16:19] = 4'd5;
    6'b010010: output_wires[16:19] = 4'd5;
    6'b010011: output_wires[16:19] = 4'd0;
    6'b010100: output_wires[16:19] = 4'd3;
    6'b010101: output_wires[16:19] = 4'd15;
    6'b010110: output_wires[16:19] = 4'd15;
    6'b010111: output_wires[16:19] = 4'd10;
    6'b011000: output_wires[16:19] = 4'd13;
    6'b011001: output_wires[16:19] = 4'd3;
    6'b011010: output_wires[16:19] = 4'd0;
    6'b011011: output_wires[16:19] = 4'd9;
    6'b011100: output_wires[16:19] = 4'd14;
    6'b011101: output_wires[16:19] = 4'd8;
    6'b011110: output_wires[16:19] = 4'd9;
    6'b011111: output_wires[16:19] = 4'd6;
    6'b100000: output_wires[16:19] = 4'd4;
    6'b100001: output_wires[16:19] = 4'd11;
    6'b100010: output_wires[16:19] = 4'd2;
    6'b100011: output_wires[16:19] = 4'd8;
    6'b100100: output_wires[16:19] = 4'd1;
    6'b100101: output_wires[16:19] = 4'd12;
    6'b100110: output_wires[16:19] = 4'd11;
    6'b100111: output_wires[16:19] = 4'd7;
    6'b101000: output_wires[16:19] = 4'd10;
    6'b101001: output_wires[16:19] = 4'd1;
    6'b101010: output_wires[16:19] = 4'd13;
    6'b101011: output_wires[16:19] = 4'd14;
    6'b101100: output_wires[16:19] = 4'd7;
    6'b101101: output_wires[16:19] = 4'd2;
    6'b101110: output_wires[16:19] = 4'd8;
    6'b101111: output_wires[16:19] = 4'd13;
    6'b110000: output_wires[16:19] = 4'd15;
    6'b110001: output_wires[16:19] = 4'd6;
    6'b110010: output_wires[16:19] = 4'd9;
    6'b110011: output_wires[16:19] = 4'd15;
    6'b110100: output_wires[16:19] = 4'd12;
    6'b110101: output_wires[16:19] = 4'd0;
    6'b110110: output_wires[16:19] = 4'd5;
    6'b110111: output_wires[16:19] = 4'd9;
    6'b111000: output_wires[16:19] = 4'd6;
    6'b111001: output_wires[16:19] = 4'd10;
    6'b111010: output_wires[16:19] = 4'd3;
    6'b111011: output_wires[16:19] = 4'd4;
    6'b111100: output_wires[16:19] = 4'd0;
    6'b111101: output_wires[16:19] = 4'd5;
    6'b111110: output_wires[16:19] = 4'd14;
    6'b111111: output_wires[16:19] = 4'd3;
endcase

case(input_wires[30:35])
    6'b000000: output_wires[20:23] = 4'd12;
    6'b000001: output_wires[20:23] = 4'd10;
    6'b000010: output_wires[20:23] = 4'd1;
    6'b000011: output_wires[20:23] = 4'd15;
    6'b000100: output_wires[20:23] = 4'd10;
    6'b000101: output_wires[20:23] = 4'd4;
    6'b000110: output_wires[20:23] = 4'd15;
    6'b000111: output_wires[20:23] = 4'd2;
    6'b001000: output_wires[20:23] = 4'd9;
    6'b001001: output_wires[20:23] = 4'd7;
    6'b001010: output_wires[20:23] = 4'd2;
    6'b001011: output_wires[20:23] = 4'd12;
    6'b001100: output_wires[20:23] = 4'd6;
    6'b001101: output_wires[20:23] = 4'd9;
    6'b001110: output_wires[20:23] = 4'd8;
    6'b001111: output_wires[20:23] = 4'd5;
    6'b010000: output_wires[20:23] = 4'd0;
    6'b010001: output_wires[20:23] = 4'd6;
    6'b010010: output_wires[20:23] = 4'd13;
    6'b010011: output_wires[20:23] = 4'd1;
    6'b010100: output_wires[20:23] = 4'd3;
    6'b010101: output_wires[20:23] = 4'd13;
    6'b010110: output_wires[20:23] = 4'd4;
    6'b010111: output_wires[20:23] = 4'd14;
    6'b011000: output_wires[20:23] = 4'd14;
    6'b011001: output_wires[20:23] = 4'd0;
    6'b011010: output_wires[20:23] = 4'd7;
    6'b011011: output_wires[20:23] = 4'd11;
    6'b011100: output_wires[20:23] = 4'd5;
    6'b011101: output_wires[20:23] = 4'd3;
    6'b011110: output_wires[20:23] = 4'd11;
    6'b011111: output_wires[20:23] = 4'd8;
    6'b100000: output_wires[20:23] = 4'd9;
    6'b100001: output_wires[20:23] = 4'd4;
    6'b100010: output_wires[20:23] = 4'd14;
    6'b100011: output_wires[20:23] = 4'd3;
    6'b100100: output_wires[20:23] = 4'd15;
    6'b100101: output_wires[20:23] = 4'd2;
    6'b100110: output_wires[20:23] = 4'd5;
    6'b100111: output_wires[20:23] = 4'd12;
    6'b101000: output_wires[20:23] = 4'd2;
    6'b101001: output_wires[20:23] = 4'd9;
    6'b101010: output_wires[20:23] = 4'd8;
    6'b101011: output_wires[20:23] = 4'd5;
    6'b101100: output_wires[20:23] = 4'd12;
    6'b101101: output_wires[20:23] = 4'd15;
    6'b101110: output_wires[20:23] = 4'd3;
    6'b101111: output_wires[20:23] = 4'd10;
    6'b110000: output_wires[20:23] = 4'd7;
    6'b110001: output_wires[20:23] = 4'd11;
    6'b110010: output_wires[20:23] = 4'd0;
    6'b110011: output_wires[20:23] = 4'd14;
    6'b110100: output_wires[20:23] = 4'd4;
    6'b110101: output_wires[20:23] = 4'd1;
    6'b110110: output_wires[20:23] = 4'd10;
    6'b110111: output_wires[20:23] = 4'd7;
    6'b111000: output_wires[20:23] = 4'd1;
    6'b111001: output_wires[20:23] = 4'd6;
    6'b111010: output_wires[20:23] = 4'd13;
    6'b111011: output_wires[20:23] = 4'd0;
    6'b111100: output_wires[20:23] = 4'd11;
    6'b111101: output_wires[20:23] = 4'd8;
    6'b111110: output_wires[20:23] = 4'd6;
    6'b111111: output_wires[20:23] = 4'd13;
endcase

case(input_wires[36:41])
    6'b000000: output_wires[24:27] = 4'd4;
    6'b000001: output_wires[24:27] = 4'd13;
    6'b000010: output_wires[24:27] = 4'd11;
    6'b000011: output_wires[24:27] = 4'd0;
    6'b000100: output_wires[24:27] = 4'd2;
    6'b000101: output_wires[24:27] = 4'd11;
    6'b000110: output_wires[24:27] = 4'd14;
    6'b000111: output_wires[24:27] = 4'd7;
    6'b001000: output_wires[24:27] = 4'd15;
    6'b001001: output_wires[24:27] = 4'd4;
    6'b001010: output_wires[24:27] = 4'd0;
    6'b001011: output_wires[24:27] = 4'd9;
    6'b001100: output_wires[24:27] = 4'd8;
    6'b001101: output_wires[24:27] = 4'd1;
    6'b001110: output_wires[24:27] = 4'd13;
    6'b001111: output_wires[24:27] = 4'd10;
    6'b010000: output_wires[24:27] = 4'd3;
    6'b010001: output_wires[24:27] = 4'd14;
    6'b010010: output_wires[24:27] = 4'd12;
    6'b010011: output_wires[24:27] = 4'd3;
    6'b010100: output_wires[24:27] = 4'd9;
    6'b010101: output_wires[24:27] = 4'd5;
    6'b010110: output_wires[24:27] = 4'd7;
    6'b010111: output_wires[24:27] = 4'd12;
    6'b011000: output_wires[24:27] = 4'd5;
    6'b011001: output_wires[24:27] = 4'd2;
    6'b011010: output_wires[24:27] = 4'd10;
    6'b011011: output_wires[24:27] = 4'd15;
    6'b011100: output_wires[24:27] = 4'd6;
    6'b011101: output_wires[24:27] = 4'd8;
    6'b011110: output_wires[24:27] = 4'd1;
    6'b011111: output_wires[24:27] = 4'd6;
    6'b100000: output_wires[24:27] = 4'd1;
    6'b100001: output_wires[24:27] = 4'd6;
    6'b100010: output_wires[24:27] = 4'd4;
    6'b100011: output_wires[24:27] = 4'd11;
    6'b100100: output_wires[24:27] = 4'd11;
    6'b100101: output_wires[24:27] = 4'd13;
    6'b100110: output_wires[24:27] = 4'd13;
    6'b100111: output_wires[24:27] = 4'd8;
    6'b101000: output_wires[24:27] = 4'd12;
    6'b101001: output_wires[24:27] = 4'd1;
    6'b101010: output_wires[24:27] = 4'd3;
    6'b101011: output_wires[24:27] = 4'd4;
    6'b101100: output_wires[24:27] = 4'd7;
    6'b101101: output_wires[24:27] = 4'd10;
    6'b101110: output_wires[24:27] = 4'd14;
    6'b101111: output_wires[24:27] = 4'd7;
    6'b110000: output_wires[24:27] = 4'd10;
    6'b110001: output_wires[24:27] = 4'd9;
    6'b110010: output_wires[24:27] = 4'd15;
    6'b110011: output_wires[24:27] = 4'd5;
    6'b110100: output_wires[24:27] = 4'd6;
    6'b110101: output_wires[24:27] = 4'd0;
    6'b110110: output_wires[24:27] = 4'd8;
    6'b110111: output_wires[24:27] = 4'd15;
    6'b111000: output_wires[24:27] = 4'd0;
    6'b111001: output_wires[24:27] = 4'd14;
    6'b111010: output_wires[24:27] = 4'd5;
    6'b111011: output_wires[24:27] = 4'd2;
    6'b111100: output_wires[24:27] = 4'd9;
    6'b111101: output_wires[24:27] = 4'd3;
    6'b111110: output_wires[24:27] = 4'd2;
    6'b111111: output_wires[24:27] = 4'd12;
endcase

case(input_wires[42:47])
    6'b000000: output_wires[28:31] = 4'd13;
    6'b000001: output_wires[28:31] = 4'd1;
    6'b000010: output_wires[28:31] = 4'd2;
    6'b000011: output_wires[28:31] = 4'd15;
    6'b000100: output_wires[28:31] = 4'd8;
    6'b000101: output_wires[28:31] = 4'd13;
    6'b000110: output_wires[28:31] = 4'd4;
    6'b000111: output_wires[28:31] = 4'd8;
    6'b001000: output_wires[28:31] = 4'd6;
    6'b001001: output_wires[28:31] = 4'd10;
    6'b001010: output_wires[28:31] = 4'd15;
    6'b001011: output_wires[28:31] = 4'd3;
    6'b001100: output_wires[28:31] = 4'd11;
    6'b001101: output_wires[28:31] = 4'd7;
    6'b001110: output_wires[28:31] = 4'd1;
    6'b001111: output_wires[28:31] = 4'd4;
    6'b010000: output_wires[28:31] = 4'd10;
    6'b010001: output_wires[28:31] = 4'd12;
    6'b010010: output_wires[28:31] = 4'd9;
    6'b010011: output_wires[28:31] = 4'd5;
    6'b010100: output_wires[28:31] = 4'd3;
    6'b010101: output_wires[28:31] = 4'd6;
    6'b010110: output_wires[28:31] = 4'd14;
    6'b010111: output_wires[28:31] = 4'd11;
    6'b011000: output_wires[28:31] = 4'd5;
    6'b011001: output_wires[28:31] = 4'd0;
    6'b011010: output_wires[28:31] = 4'd0;
    6'b011011: output_wires[28:31] = 4'd14;
    6'b011100: output_wires[28:31] = 4'd12;
    6'b011101: output_wires[28:31] = 4'd9;
    6'b011110: output_wires[28:31] = 4'd7;
    6'b011111: output_wires[28:31] = 4'd2;
    6'b100000: output_wires[28:31] = 4'd7;
    6'b100001: output_wires[28:31] = 4'd2;
    6'b100010: output_wires[28:31] = 4'd11;
    6'b100011: output_wires[28:31] = 4'd1;
    6'b100100: output_wires[28:31] = 4'd4;
    6'b100101: output_wires[28:31] = 4'd14;
    6'b100110: output_wires[28:31] = 4'd1;
    6'b100111: output_wires[28:31] = 4'd7;
    6'b101000: output_wires[28:31] = 4'd9;
    6'b101001: output_wires[28:31] = 4'd4;
    6'b101010: output_wires[28:31] = 4'd12;
    6'b101011: output_wires[28:31] = 4'd10;
    6'b101100: output_wires[28:31] = 4'd14;
    6'b101101: output_wires[28:31] = 4'd8;
    6'b101110: output_wires[28:31] = 4'd2;
    6'b101111: output_wires[28:31] = 4'd13;
    6'b110000: output_wires[28:31] = 4'd0;
    6'b110001: output_wires[28:31] = 4'd15;
    6'b110010: output_wires[28:31] = 4'd6;
    6'b110011: output_wires[28:31] = 4'd12;
    6'b110100: output_wires[28:31] = 4'd10;
    6'b110101: output_wires[28:31] = 4'd9;
    6'b110110: output_wires[28:31] = 4'd13;
    6'b110111: output_wires[28:31] = 4'd0;
    6'b111000: output_wires[28:31] = 4'd15;
    6'b111001: output_wires[28:31] = 4'd3;
    6'b111010: output_wires[28:31] = 4'd3;
    6'b111011: output_wires[28:31] = 4'd5;
    6'b111100: output_wires[28:31] = 4'd5;
    6'b111101: output_wires[28:31] = 4'd6;
    6'b111110: output_wires[28:31] = 4'd8;
    6'b111111: output_wires[28:31] = 4'd11;
endcase


end

endmodule
