// $Id: $
// File name:   tb_control.sv
// Created:     4/12/2015
// Author:      Lucas Dahl
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: tb for controller

`timescale 1ns / 100ps

module tb_control();

	parameter CLK_PERIOD = 2.5;

	reg tb_clk;
	reg tb_n_rst;
	reg [63:0] tb_data_in;
	reg tb_start;
	reg [63:0] tb_data_out;
	reg [2:0] tb_mode;
	reg tb_data_ready;
	reg tb_estart;
	reg tb_edone;
	reg [163:0] tb_k;
	reg [163:0] tb_Pix;
	reg [163:0] tb_Piy;
	reg [163:0] tb_Pox;
	reg [163:0] tb_Poy;
	reg [63:0] tb_DES_output;
	reg [63:0] tb_DES_input;
	reg [163:0] tb_Skx;
	reg [163:0] tb_Sky;

	
	control DUT(.clk(tb_clk), .n_rst(tb_n_rst), .start(tb_start), .data_in(tb_data_in), .mode(tb_mode), .data_out(tb_data_out), .data_ready(tb_data_ready), .edone(tb_edone), .Pox(tb_Pox), .Poy(tb_Poy), .k(tb_k), .Pix(tb_Pix), .Piy(tb_Piy), .estart(tb_estart), .DES_output(tb_DES_output), .Skx(tb_Skx), .Sky(tb_Sky), .DES_input(tb_DES_input));

	always
	begin : CLK_GEN
		tb_clk = 1'b0;
		#(CLK_PERIOD / 2);
		tb_clk = 1'b1;
		#(CLK_PERIOD / 2);
	end


	initial
	begin
		tb_edone = 1'b1;
		tb_n_rst = 1'b0;
		#CLK_PERIOD;
		#CLK_PERIOD;
		tb_n_rst = 1'b1;
		tb_start = 1'b0;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1010101010101010101010101010101010101010101010101010101010101010;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		tb_edone = 1'b1;
		#CLK_PERIOD;
		tb_edone = 1'b0;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		tb_start = 1'b1;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1111111111111111111111111111111111111111111111111111111111111111;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		#CLK_PERIOD;
		tb_data_in = 64'b1010101010101010101010101010101010101010101010101010101010101010;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		tb_edone = 1'b1;
		#CLK_PERIOD;
		tb_edone = 1'b0;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		tb_data_in = 64'b1100110101111010101010101010101010101010100101011001010010101010;
		#CLK_PERIOD;
		tb_data_in = 64'b1010101010101010101010110101001110101011101000000000101010101010;
		#CLK_PERIOD;
		tb_data_in = 64'b0000000000000000000000000000000000000000101010101010101010101010;
		#CLK_PERIOD;
		tb_data_in = 64'b1010101111111111111111111111111111111111111110000000001010101010;
		#CLK_PERIOD;
		tb_data_in = 64'b1010101010101010101011111111111010101010101010101010101010101010;
		#CLK_PERIOD;
		tb_data_in = 64'b1010100010101011011111101010101010101010101010101010100000101010;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		#CLK_PERIOD;
		tb_start = 1'b0;
		#CLK_PERIOD;
		#CLK_PERIOD;
		
	end
endmodule
